`timescale 1ns / 1ps
//This is a tempplate from the instructor
//HUST Fall 2020
//Read==1
//Write==0
module I2C_SDAmodule(input ReadorWrite, Select, StartStopAck, ShiftOut,
output ShiftIn, inout SDA);



	
endmodule
